module sending_tx(
    input wire clk,
    input wire [31:0] xo,
    input wire [31:0] xt,
    input wire [31:0] yo,
    input wire [31:0] yt,
    input wire g_send,
    input wire [1:0] intensity,
    input wire reset,
    input wire BTNU,
    input wire BTNL,
    input wire BTNR,
    input wire BTND,
    input wire rx,
    output wire tx,
    output wire busy
);
    assign busy = g_busy || uart_tx_busy;
    wire uart_tx_busy;
    wire tx_valid, button_valid, g_valid;

    wire g_busy, b_busy, ready_send;

    wire[7:0] test_letter, g_letter, b_letter, rx_data;
    
    assign tx_valid = (g_busy) ? g_valid : b_valid;
    assign test_letter = (g_busy) ? g_letter : b_letter;
    
    button_send sending_button(
        .clk(clk),
        .reset(reset),
        .BTNU(BTNU), 
        .BTNL(BTNL),
        .BTNR(BTNR),
        .BTND(BTND),
        .tx_ready(!uart_tx_busy && !g_busy),
        .tx_valid(b_valid),
        .tx_data(b_letter)
);

    uart_receive urt(
        .clk(clk),
        .reset(reset),
        .rx(rx),
        .rx_done(rx_done),
        .rx_data(rx_data)
    );

    check_receive okay(
        .clk(clk),
        .reset(reset),
        .rx_data(rx_data),
        .rx_done(rx_done),
        .ready_send(ready_send)
    );

    uart_transmit uut(
        .clk(clk), 
        .reset(reset), 
        .tx_send(tx), 
        .tx_busy(uart_tx_busy), 
        .tx_start(tx_valid), 
        .tx_data(test_letter));

    gcode_sender getting_gcode(
        .xo(xo),
        .xt(xt),
        .yo(yo),
        .yt(yt),
        .intensity(intensity),
        .receive_ok(1'b1),
        .g_send(g_send),
        .g_busy(g_busy),
        .clk(clk),
        .reset(reset),
        .tx_ready(!uart_tx_busy),
        .tx_valid(g_valid),
        .tx_data(g_letter));
endmodule