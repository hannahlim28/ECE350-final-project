module or32(output [31:0] y, input [31:0] a, input [31:0] b);  
  or  ORbit[31:0](y, a, b);

endmodule