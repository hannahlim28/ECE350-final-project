module not32(output [31:0] y, input [31:0] a);
  not NOTbit[31:0](y, a);

endmodule
